library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library unisim;
use unisim.vcomponents.all;
use work.miningshell_types.all;


-- This unit wraps a pair of MMCMs and a BUFGMUX to allow for seamless adjustment
-- of clocks used by the hashing core. It basically has the capabilities of one MMCM,
-- i.e. it could have up to 6 clock outputs with different capabilities. It works
-- by reconfiguring the currently unused MMCM while the hashing core is running on
-- clocks generated by the other one, waiting for the reconfigured MCMM to lock,
-- and then switching the clock outputs over to the reconfigured MMCM using the
-- BUFGMUX, so that the other MMCM can be reconfigured for the next adjustment.
-- The DRP signals for reconfiguration and the multiplexer control signal are
-- provided by the shell and are just routed to the MMCMs by this module.
-- This reference implementation only uses the first output of the MMCM,
-- but adding further output channels is quite straightforward.
entity clkgen is
  port(
    refclk : in std_logic;  -- Reference clock for MMCMs
    to_clkgen : in to_clkgen;  -- MMCM/MUX control signals from the shell
    from_clkgen : out from_clkgen;  -- MMCM status signals to the shell
    hashing_clk : out std_Logic  -- Output clock (hashing core clock)
  );
end clkgen;


architecture structure of clkgen is

  -- Output signals of the first MMCM
  signal mmcm0_fb : std_logic;
  signal mmcm0_out0 : std_logic;

  -- Output signals of the second MMCM
  signal mmcm1_fb : std_logic;
  signal mmcm1_out0 : std_logic;

begin

  -- First MMCM (the generic values are just set to make synthesis happy, the MMCM
  -- will be reconfigured by software before being started for the first time)
  mmcm0 : MMCME4_ADV
    generic map (
      CLKIN1_PERIOD => 3.333,
      DIVCLK_DIVIDE => 3,
      CLKFBOUT_MULT_F => 10.0,
      CLKOUT0_DIVIDE_F => 5.0
    )
    port map (
      RST => to_clkgen.pll_drp(0).rst,
      PWRDWN => to_clkgen.pll_drp(0).pwrdwn,
      CLKIN1 => refclk,
      CLKIN2 => '0',
      CLKINSEL => '1',
      CLKFBOUT => mmcm0_fb,
      CLKFBIN => mmcm0_fb,
      CLKFBOUTB => open,
      CLKFBSTOPPED => open,
      CLKINSTOPPED => open,
      LOCKED => from_clkgen.pll_drp(0).locked,
      CLKOUT0 => mmcm0_out0,
      CLKOUT0B => open,
      CLKOUT1 => open,
      CLKOUT1B => open,
      CLKOUT2 => open,
      CLKOUT2B => open,
      CLKOUT3 => open,
      CLKOUT3B => open,
      CLKOUT4 => open,
      CLKOUT5 => open,
      CLKOUT6 => open,
      DCLK => to_clkgen.pll_drp(0).dclk,
      DRDY => from_clkgen.pll_drp(0).drdy,
      DEN => to_clkgen.pll_drp(0).den,
      DWE => to_clkgen.pll_drp(0).dwe,
      DADDR => to_clkgen.pll_drp(0).daddr,
      DI => to_clkgen.pll_drp(0).di,
      DO => from_clkgen.pll_drp(0).do,
      PSDONE => open,
      PSCLK => '0',
      PSEN => '0',
      PSINCDEC => '0',
      CDDCDONE => open,
      CDDCREQ => '0'
    );

  -- Second MMCM (the generic values are just set to make synthesis happy, the MMCM
  -- will be reconfigured by software before being started for the first time)
  mmcm1 : MMCME4_ADV
    generic map (
      CLKIN1_PERIOD => 3.333,
      DIVCLK_DIVIDE => 3,
      CLKFBOUT_MULT_F => 10.0,
      CLKOUT0_DIVIDE_F => 5.0
    )
    port map (
      RST => to_clkgen.pll_drp(1).rst,
      PWRDWN => to_clkgen.pll_drp(1).pwrdwn,
      CLKIN1 => refclk,
      CLKIN2 => '0',
      CLKINSEL => '1',
      CLKFBOUT => mmcm1_fb,
      CLKFBIN => mmcm1_fb,
      CLKFBOUTB => open,
      CLKFBSTOPPED => open,
      CLKINSTOPPED => open,
      LOCKED => from_clkgen.pll_drp(1).locked,
      CLKOUT0 => mmcm1_out0,
      CLKOUT0B => open,
      CLKOUT1 => open,
      CLKOUT1B => open,
      CLKOUT2 => open,
      CLKOUT2B => open,
      CLKOUT3 => open,
      CLKOUT3B => open,
      CLKOUT4 => open,
      CLKOUT5 => open,
      CLKOUT6 => open,
      DCLK => to_clkgen.pll_drp(1).dclk,
      DRDY => from_clkgen.pll_drp(1).drdy,
      DEN => to_clkgen.pll_drp(1).den,
      DWE => to_clkgen.pll_drp(1).dwe,
      DADDR => to_clkgen.pll_drp(1).daddr,
      DI => to_clkgen.pll_drp(1).di,
      DO => from_clkgen.pll_drp(1).do,
      PSDONE => open,
      PSCLK => '0',
      PSEN => '0',
      PSINCDEC => '0',
      CDDCDONE => open,
      CDDCREQ => '0'
    );

  -- Multiplexer for the first (and only) output channel (add more as needed)
  mmcm_mux : BUFGMUX port map(I0 => mmcm0_out0, I1 => mmcm1_out0, S => to_clkgen.mux_sel, O => hashing_clk);

end structure;
